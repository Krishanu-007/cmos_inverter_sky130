.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.include /home/krishanu/Desktop/cmos_inverter_sky130/Simulation/Layout_Simulations/inv_layout_fixed.spice
Vdd Vdd 0 1.8
Vin Vin 0 0
Xinv Vin Vout Vdd 0 inv_layout_fixed
Cload Vout 0 10f
.dc Vin 0 1.8 1m
.save all
.end

