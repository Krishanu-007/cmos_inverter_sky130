** sch_path: /home/krish/Desktop/cmos_inverter_sky130/Xschem/power.sch
**.subckt power
x1 Vdd Vin Vout GND inv
Vdd Vdd GND 1.8
Vin Vin GND PULSE(0 1.8 0 500ps 500ps 4ns 10ns)
C1 Vout GND 100f m=1
**** begin user architecture code

.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.tran 100ps 30ns
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/krish/Desktop/cmos_inverter_sky130/Xschem/inv.sym
** sch_path: /home/krish/Desktop/cmos_inverter_sky130/Xschem/inv.sch
.subckt inv Vdd Vin Vout Vss
*.ipin Vin
*.ipin Vss
*.ipin Vdd
*.opin Vout
XM1 Vout Vin Vss GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin Vdd VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
